library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

 
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI  : std_logic_vector(3 downto 0) := "0100";
  constant STA  : std_logic_vector(3 downto 0) := "0101";
  constant JMP  : std_logic_vector(3 downto 0) := "0110";
  constant JEQ  : std_logic_vector(3 downto 0) := "0111";
  constant CEQ  : std_logic_vector(3 downto 0) := "1000";
  constant JSR  : std_logic_vector(3 downto 0) := "1001";
  constant RET  : std_logic_vector(3 downto 0) := "1010";
   constant OP_AND:std_logic_vector(3 downto 0) := "1011";


  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
-- RESET:
tmp(1) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(2) := x"5" & "00" & '0'& '1' & x"FE";	-- STA @510 	# Limpando key 1
tmp(3) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando segundos
tmp(4) := x"5" & "00" & '0'& '0' & x"00";	-- STA @0 	# Limpando endereço de unidade
tmp(5) := x"5" & "00" & '0'& '0' & x"01";	-- STA @1 	# Limpando endereço de dezena
tmp(6) := x"5" & "00" & '0'& '0' & x"02";	-- STA @2 	# Limpando endereço de centena
tmp(7) := x"5" & "00" & '0'& '0' & x"03";	-- STA @3 	# Limpando endereço de milhar
tmp(8) := x"5" & "00" & '0'& '0' & x"04";	-- STA @4 	# Limpando endereço de dezena de milhar
tmp(9) := x"5" & "00" & '0'& '0' & x"05";	-- STA @5 	# Limpando endereço de centena de milhar
tmp(10) := x"5" & "00" & '0'& '1' & x"20";	-- STA @288 	# Limpando endereço do HEX0
tmp(11) := x"5" & "00" & '0'& '1' & x"21";	-- STA @289 	# Limpando endereço do HEX1
tmp(12) := x"5" & "00" & '0'& '1' & x"22";	-- STA @290 	# Limpando endereço do HEX2
tmp(13) := x"5" & "00" & '0'& '1' & x"23";	-- STA @291 	# Limpando endereço do HEX3
tmp(14) := x"5" & "00" & '0'& '1' & x"24";	-- STA @292 	# Limpando endereço do HEX4
tmp(15) := x"5" & "00" & '0'& '1' & x"25";	-- STA @293 	# Limpando endereço do HEX5
tmp(16) := x"5" & "00" & '1' & '1' & x"FF";	-- STA @1023 	# Limpando endereço do BUZZER
tmp(17) := x"4" & "00" & '0'& '0' & x"07";	-- LDI $7 	# Carregando 7 no acumulador
tmp(18) := x"5" & "00" & '0'& '0' & x"84";	-- STA @132 	# Liga cor
tmp(19) := x"4" & "00" & '0'& '0' & x"05";	-- LDI $5 	# Carregando 3 no acumulador
tmp(20) := x"5" & "00" & '0'& '0' & x"80";	-- STA @128 	# Carregando 3 na LINHA
tmp(21) := x"4" & "00" & '0'& '0' & x"0B";	-- LDI $11 	# Carregando 9 no acumulador
tmp(22) := x"5" & "00" & '0'& '0' & x"81";	-- STA @129 	# Carregando 9 na COLUNA
tmp(23) := x"4" & "00" & '0'& '0' & x"1A";	-- LDI $26 	# Carregando : no acumulador
tmp(24) := x"5" & "00" & '0'& '0' & x"82";	-- STA @130 	# Carregando : na posição 130
tmp(25) := x"5" & "00" & '0'& '0' & x"83";	-- STA @131 	# Liga VGA
tmp(26) := x"4" & "00" & '0'& '0' & x"08";	-- LDI $8 	# Carregando 9 no acumulador
tmp(27) := x"5" & "00" & '0'& '0' & x"81";	-- STA @129 	# Carregando 9 na COLUNA
tmp(28) := x"4" & "00" & '0'& '0' & x"1A";	-- LDI $26 	# Carregando : no acumulador
tmp(29) := x"5" & "00" & '0'& '0' & x"82";	-- STA @130 	# Carregando : na posição 130
tmp(30) := x"5" & "00" & '0'& '0' & x"83";	-- STA @131 	# Liga VGA
tmp(31) := x"4" & "00" & '0'& '0' & x"02";	-- LDI $2 	# Carregando 2 no acumulador
tmp(32) := x"5" & "00" & '0'& '0' & x"34";	-- STA @52 	# Carregando 2 na posição 52
tmp(33) := x"4" & "00" & '0'& '0' & x"03";	-- LDI $3 	# Carregando 4 no acumulador
tmp(34) := x"5" & "00" & '0'& '0' & x"35";	-- STA @53 	# Carregando 4 na posição 53
tmp(35) := x"4" & "00" & '0'& '0' & x"04";	-- LDI $4 	# Carregando 4 no acumulador
tmp(36) := x"5" & "00" & '0'& '0' & x"36";	-- STA @54 	# Carregando 4 na posição 54
tmp(37) := x"4" & "00" & '0'& '0' & x"05";	-- LDI $5 	# Carregando 5 no acumulador
tmp(38) := x"5" & "00" & '0'& '0' & x"37";	-- STA @55 	# Carregando 5 na posição 55
tmp(39) := x"4" & "00" & '0'& '0' & x"09";	-- LDI $9 	# Carregando 9 no acumulador
tmp(40) := x"5" & "00" & '0'& '0' & x"3B";	-- STA @59 	# Carregando 9 na posição 59
tmp(41) := x"4" & "00" & '0'& '0' & x"0A";	-- LDI $10 	# Carregando 10 no acumulador
tmp(42) := x"5" & "00" & '0'& '0' & x"3C";	-- STA @60 	# Carergando 10 na posição 60
tmp(43) := x"4" & "00" & '0'& '0' & x"01";	-- LDI $1 	# Carregando 1 no acumulador
tmp(44) := x"5" & "00" & '0'& '0' & x"33";	-- STA @51 	# Carregando 1 na posição 51
tmp(45) := x"4" & "00" & '0'& '0' & x"09";	-- LDI $9
tmp(46) := x"5" & "00" & '0'& '0' & x"28";	-- STA @40 	# Limpando endereço de temp 1
tmp(47) := x"5" & "00" & '0'& '0' & x"0A";	-- STA @10 	# Limite das unidades
tmp(48) := x"5" & "00" & '0'& '0' & x"0C";	-- STA @12 	# Limite das centenas
tmp(49) := x"5" & "00" & '0'& '0' & x"2A";	-- STA @42 	# Limpando endereço de temp 3
tmp(50) := x"4" & "00" & '0'& '0' & x"05";	-- LDI $5 
tmp(51) := x"5" & "00" & '0'& '0' & x"0B";	-- STA @11 	# Limite das dezenas
tmp(52) := x"5" & "00" & '0'& '0' & x"29";	-- STA @41 	# Limpando endereço de temp 2
tmp(53) := x"5" & "00" & '0'& '0' & x"0D";	-- STA @13 	# Limite dos milhares
tmp(54) := x"5" & "00" & '0'& '0' & x"2B";	-- STA @43 	# Limpando endereço de temp 4
tmp(55) := x"4" & "00" & '0'& '0' & x"03";	-- LDI $3 
tmp(56) := x"5" & "00" & '0'& '0' & x"0E";	-- STA @14 	# Limite das dezenas de milhares
tmp(57) := x"5" & "00" & '0'& '0' & x"2C";	-- STA @44 	# Limpando endereço de temp 5
tmp(58) := x"4" & "00" & '0'& '0' & x"02";	-- LDI $2
tmp(59) := x"5" & "00" & '0'& '0' & x"0F";	-- STA @15 	# Limite das centenas de milhares
tmp(60) := x"5" & "00" & '0'& '0' & x"2D";	-- STA @45 	# Limpando endereço de temp 6
tmp(61) := x"4" & "00" & '0'& '0' & x"63";	-- LDI $99 	# Carregando 99 no acumulador
tmp(62) := x"5" & "00" & '0'& '0' & x"1D";	-- STA @29 	# Carregando 100 na posição 29
tmp(63) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carregando 0 no acumulador
tmp(64) := x"5" & "00" & '0'& '1' & x"F4";	-- STA @500 	# Desligando o display 0
tmp(65) := x"5" & "00" & '0'& '0' & x"14";	-- STA @20 	#temporizador 1
tmp(66) := x"5" & "00" & '0'& '0' & x"15";	-- STA @21 	#temporizador 2
tmp(67) := x"5" & "00" & '0'& '0' & x"16";	-- STA @22 	#temporizador 3
tmp(68) := x"5" & "00" & '0'& '0' & x"17";	-- STA @23 	# PISCA OU NÃO PISCA
tmp(69) := x"6" & "00"& '0' & '1' & x"7D";	-- JMP %le_key 	# Vai para o label le_key
-- temporizador_1_segundo:
tmp(71) := x"1" & "00" & '0'& '0' & x"14";	-- LDA @20 	# Carrega o acumulador com o endereço de temporizador 1
tmp(72) := x"8" & "00" & '0'& '0' & x"1D";	-- CEQ @29 	# Compara o valor do acumulador com o valor 99
tmp(73) := x"7" & "00" & '0' & '0' & x"4E";	-- JEQ %temporizador_2_segundo 	# Se for igual, vai para o label temporizador_2_segundo
tmp(74) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(75) := x"5" & "00" & '0'& '0' & x"14";	-- STA @20 	# Armazena o valor do acumulador no endereço de temporizador 1
tmp(76) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- temporizador_2_segundo:
tmp(78) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(79) := x"5" & "00" & '0'& '0' & x"14";	-- STA @20 	# Armazena o valor do acumulador no endereço de temporizador 1
tmp(80) := x"1" & "00" & '0'& '0' & x"15";	-- LDA @21 	# Carrega o acumulador com o endereço de temporizador 2
tmp(81) := x"8" & "00" & '0'& '0' & x"1D";	-- CEQ @29 	# Compara o valor do acumulador com o valor 99
tmp(82) := x"7" & "00" & '0' & '0' & x"57";	-- JEQ %temporizador_3_segundo 	# Se for igual, vai para o label temporizador_3_segundo
tmp(83) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(84) := x"5" & "00" & '0'& '0' & x"15";	-- STA @21 	# Armazena o valor do acumulador no endereço de temporizador 2
tmp(85) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- temporizador_3_segundo:
tmp(87) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(88) := x"5" & "00" & '0'& '0' & x"15";	-- STA @21 	# Armazena o valor do acumulador no endereço de temporizador 2
tmp(89) := x"1" & "00" & '0'& '0' & x"16";	-- LDA @22 	# Carrega o acumulador com o endereço de temporizador 3
tmp(90) := x"8" & "00" & '0'& '0' & x"1D";	-- CEQ @29 	# Compara o valor do acumulador com o valor 99
tmp(91) := x"7" & "00" & '0' & '0' & x"60";	-- JEQ %PISCA 	# Se for igual, vai para o label LIMPA
tmp(92) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(93) := x"5" & "00" & '0'& '0' & x"16";	-- STA @22 	# Armazena o valor do acumulador no endereço de temporizador 3
tmp(94) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- PISCA:
tmp(96) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(97) := x"5" & "00" & '0'& '0' & x"16";	-- STA @22 	# Limpando temporizador 3
tmp(98) := x"1" & "00" & '0'& '0' & x"17";	-- LDA @23 	# Carrega o acumulador com o endereço de PISCA
tmp(99) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(100) := x"7" & "00" & '0' & '0' & x"69";	-- JEQ %LIMPA 	# Se for igual, vai para o label LIMPA
tmp(101) := x"4" & "00" & '0'& '0' & x"01";	-- LDI $1 	# Carrega 1 no acumulador
tmp(102) := x"5" & "00" & '0'& '0' & x"17";	-- STA @23 	# Armazena o valor do acumulador no endereço de PISCA
tmp(103) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- LIMPA:
tmp(105) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(106) := x"5" & "00" & '0'& '0' & x"17";	-- STA @23 	# Armazena o valor do acumulador no endereço de PISCA
tmp(107) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- define_limites_unidades:
tmp(109) := x"5" & "00" & '0'& '1' & x"FE";	-- STA @510 	# Limpando key 1
tmp(110) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(111) := x"9" & "00" & '1' & '0' & x"6E";	-- JSR %atualiza_displays_limites 	# Vai para o label atualiza_displays_limites
-- checa_limites_unidades:
tmp(113) := x"9" & "00" & '0' & '0' & x"47";	-- JSR %temporizador_1_segundo 	# Vai para o label temporizador_1_segundo
tmp(114) := x"1" & "00" & '0'& '0' & x"17";	-- LDA @23 	# Carrega o acumulador com o endereço de PISCA
tmp(115) := x"5" & "00" & '0'& '1' & x"F4";	-- STA @500 	# Desliga o display unidade
tmp(116) := x"1" & "00" & '0'& '1' & x"61";	-- LDA @353 	# Carrega o acumulador com o key 1
tmp(117) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(118) := x"7" & "00" & '0' & '0' & x"89";	-- JEQ %define_limites_dezenas 	# Se for igual, vai para o label define_limites_dezenas
tmp(119) := x"1" & "00" & '0'& '1' & x"60";	-- LDA @352 	# Carrega o acumulador com o key 0
tmp(120) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador com o valor 0
tmp(121) := x"7" & "00" & '0' & '0' & x"71";	-- JEQ %checa_limites_unidades 	# Se for igual, vai para o label checa_limites_unidades
tmp(122) := x"9" & "00" & '0' & '0' & x"7D";	-- JSR %adiciona_unidade 	# Se não for igual, vai para o label adiciona_unidade
tmp(123) := x"6" & "00" & '0' & '0' & x"6D";	-- JMP %define_limites_unidades 	# Se não for igual, volta para o label define_limites_unidades
-- adiciona_unidade:
tmp(125) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(126) := x"1" & "00" & '0'& '0' & x"28";	-- LDA @40 	# Carrega o acumulador com o endereço de Limite de unidade
tmp(127) := x"8" & "00" & '0'& '0' & x"3B";	-- CEQ @59 	# Compara o valor do acumulador com o valor 9
tmp(128) := x"7" & "00" & '0' & '0' & x"85";	-- JEQ %zera_unidade 	# Se for igual, vai para o label zera_unidade
tmp(129) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(130) := x"5" & "00" & '0'& '0' & x"28";	-- STA @40 	# Armazena o valor do acumulador no endereço de Limite de unidade
tmp(131) := x"A" & "00" & '0' & '0' & x"00";	-- RET 
-- zera_unidade:
tmp(133) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(134) := x"5" & "00" & '0'& '0' & x"28";	-- STA @40 	# Armazena o valor do acumulador no endereço de Limite de unidade
tmp(135) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- define_limites_dezenas:
tmp(137) := x"5" & "00" & '0'& '1' & x"FE";	-- STA @510 	# Limpando key 1
tmp(138) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(139) := x"9" & "00" & '1' & '0' & x"6E";	-- JSR %atualiza_displays_limites 	# Vai para o label atualiza_displays_limites
-- checa_limites_dezenas:
tmp(141) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(142) := x"5" & "00" & '0'& '1' & x"F4";	-- STA @500 	# liga o display unidade
tmp(143) := x"9" & "00" & '0' & '0' & x"47";	-- JSR %temporizador_1_segundo 	# Vai para o label temporizador_1_segundo
tmp(144) := x"1" & "00" & '0'& '0' & x"17";	-- LDA @23 	# Carrega o acumulador com o endereço de PISCA
tmp(145) := x"5" & "00" & '0'& '1' & x"F5";	-- STA @501 	# Desliga o display unidade
tmp(146) := x"1" & "00" & '0'& '1' & x"61";	-- LDA @353 	# Carrega o acumulador com o key 1
tmp(147) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(148) := x"7" & "00" & '0' & '0' & x"A6";	-- JEQ %define_limites_centenas 	# Se for igual, vai para o label define_limites_dezenas
tmp(149) := x"1" & "00" & '0'& '1' & x"60";	-- LDA @352 	# Carrega o acumulador com o key 0
tmp(150) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador com o valor 0
tmp(151) := x"7" & "00" & '0' & '0' & x"8D";	-- JEQ %checa_limites_dezenas 	# Se for igual, vai para o label checa_limites_dezenas
tmp(152) := x"9" & "00" & '0' & '0' & x"9C";	-- JSR %adiciona_dezena 	# Se não for igual, vai para o label adiciona_dezena
tmp(153) := x"5" & "00" & '0'& '0' & x"29";	-- STA @41 	# Armazena o valor do acumulador no endereço de Limite de dezenas
tmp(154) := x"6" & "00" & '0' & '0' & x"89";	-- JMP %define_limites_dezenas 	# Se não for igual, volta para o label define_limites_dezenas
-- adiciona_dezena:
tmp(156) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(157) := x"1" & "00" & '0'& '0' & x"29";	-- LDA @41 	# Carrega o acumulador com o endereço de Limite de dezena
tmp(158) := x"8" & "00" & '0'& '0' & x"37";	-- CEQ @55 	# Compara o valor do acumulador com o valor 5
tmp(159) := x"7" & "00" & '0' & '0' & x"A3";	-- JEQ %zera_dezena 	# Se for igual, vai para o label zera_dezena
tmp(160) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(161) := x"A" & "00" & '0' & '0' & x"00";	-- RET 
-- zera_dezena:
tmp(163) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(164) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- define_limites_centenas:
tmp(166) := x"5" & "00" & '0'& '1' & x"FE";	-- STA @510 	# Limpando key 1
tmp(167) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(168) := x"9" & "00" & '1' & '0' & x"6E";	-- JSR %atualiza_displays_limites 	# Vai para o label atualiza_displays_limites
-- checa_limites_centenas:
tmp(170) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(171) := x"5" & "00" & '0'& '1' & x"F5";	-- STA @501 	# liga o display DEZENA
tmp(172) := x"9" & "00" & '0' & '0' & x"47";	-- JSR %temporizador_1_segundo 	# Vai para o label temporizador_1_segundo
tmp(173) := x"1" & "00" & '0'& '0' & x"17";	-- LDA @23 	# Carrega o acumulador com o endereço de PISCA
tmp(174) := x"5" & "00" & '0'& '1' & x"F6";	-- STA @502 	# Desliga o display unidade
tmp(175) := x"1" & "00" & '0'& '1' & x"61";	-- LDA @353 	# Carrega o acumulador com o key 1
tmp(176) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(177) := x"7" & "00" & '0' & '0' & x"C3";	-- JEQ %define_limites_milhares 	# Se for igual, vai para o label define_limites_centenas
tmp(178) := x"1" & "00" & '0'& '1' & x"60";	-- LDA @352 	# Carrega o acumulador com o key 0
tmp(179) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador com o valor 0
tmp(180) := x"7" & "00" & '0' & '0' & x"AA";	-- JEQ %checa_limites_centenas 	# Se for igual, vai para o label checa_limites_centenas
tmp(181) := x"9" & "00" & '0' & '0' & x"B9";	-- JSR %adiciona_centena 	# Se não for igual, vai para o label adiciona_centena
tmp(182) := x"5" & "00" & '0'& '0' & x"2A";	-- STA @42 	# Armazena o valor do acumulador no endereço de Limite de centenas
tmp(183) := x"6" & "00" & '0' & '0' & x"A6";	-- JMP %define_limites_centenas 	# Se não for igual, volta para o label define_limites_centenas
-- adiciona_centena:
tmp(185) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(186) := x"1" & "00" & '0'& '0' & x"2A";	-- LDA @42 	# Carrega o acumulador com o endereço de Limite de centena
tmp(187) := x"8" & "00" & '0'& '0' & x"3B";	-- CEQ @59 	# Compara o valor do acumulador com o valor 9
tmp(188) := x"7" & "00" & '0' & '0' & x"C0";	-- JEQ %zera_centena 	# Se for igual, vai para o label zera_centena
tmp(189) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(190) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- zera_centena:
tmp(192) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(193) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- define_limites_milhares:
tmp(195) := x"5" & "00" & '0'& '1' & x"FE";	-- STA @510 	# Limpando key 1
tmp(196) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(197) := x"9" & "00" & '1' & '0' & x"6E";	-- JSR %atualiza_displays_limites 	# Vai para o label atualiza_displays_limites
-- checa_limites_milhares:
tmp(199) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(200) := x"5" & "00" & '0'& '1' & x"F6";	-- STA @502 	# liga o display unidade
tmp(201) := x"9" & "00" & '0' & '0' & x"47";	-- JSR %temporizador_1_segundo 	# Vai para o label temporizador_1_segundo
tmp(202) := x"1" & "00" & '0'& '0' & x"17";	-- LDA @23 	# Carrega o acumulador com o endereço de PISCA
tmp(203) := x"5" & "00" & '0'& '1' & x"F7";	-- STA @503 	# Desliga o display unidade
tmp(204) := x"1" & "00" & '0'& '1' & x"61";	-- LDA @353 	# Carrega o acumulador com o key 1
tmp(205) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(206) := x"7" & "00" & '0' & '0' & x"E0";	-- JEQ %define_limites_dezenas_de_milhares 	# Se for igual, vai para o label define_limites_milhares
tmp(207) := x"1" & "00" & '0'& '1' & x"60";	-- LDA @352 	# Carrega o acumulador com o key 0
tmp(208) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador com o valor 0
tmp(209) := x"7" & "00" & '0' & '0' & x"C7";	-- JEQ %checa_limites_milhares 	# Se for igual, vai para o label checa_limites_milhares
tmp(210) := x"9" & "00" & '0' & '0' & x"D6";	-- JSR %adiciona_milhar 	# Se não for igual, vai para o label adiciona_milhar
tmp(211) := x"5" & "00" & '0'& '0' & x"2B";	-- STA @43 	# Armazena o valor do acumulador no endereço de Limite de milhares
tmp(212) := x"6" & "00" & '0' & '0' & x"C3";	-- JMP %define_limites_milhares 	# Se não for igual, volta para o label define_limites_milhares
-- adiciona_milhar:
tmp(214) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(215) := x"1" & "00" & '0'& '0' & x"2B";	-- LDA @43 	# Carrega o acumulador com o endereço de Limite de milhar
tmp(216) := x"8" & "00" & '0'& '0' & x"37";	-- CEQ @55 	# Compara o valor do acumulador com o valor 9
tmp(217) := x"7" & "00" & '0' & '0' & x"DD";	-- JEQ %zera_milhar 	# Se for igual, vai para o label zera_milhar
tmp(218) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(219) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- zera_milhar:
tmp(221) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(222) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- define_limites_dezenas_de_milhares:
tmp(224) := x"5" & "00" & '0'& '1' & x"FE";	-- STA @510 	# Limpando key 1
tmp(225) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(226) := x"9" & "00" & '1' & '0' & x"6E";	-- JSR %atualiza_displays_limites 	# Vai para o label atualiza_displays_limites
-- checa_limites_dezenas_de_milhares:
tmp(228) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(229) := x"5" & "00" & '0'& '1' & x"F7";	-- STA @503 	# liga o display unidade
tmp(230) := x"9" & "00" & '0' & '0' & x"47";	-- JSR %temporizador_1_segundo 	# Vai para o label temporizador_1_segundo
tmp(231) := x"1" & "00" & '0'& '0' & x"17";	-- LDA @23 	# Carrega o acumulador com o endereço de PISCA
tmp(232) := x"5" & "00" & '0'& '1' & x"F8";	-- STA @504 	# Desliga o display unidade
tmp(233) := x"1" & "00" & '0'& '1' & x"61";	-- LDA @353 	# Carrega o acumulador com o key 1
tmp(234) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(235) := x"7" & "00"& '0' & '1' & x"06";	-- JEQ %define_limites_centenas_de_milhares 	# Se for igual, vai para o label define_limites_dezenas_de_milhares
tmp(236) := x"1" & "00" & '0'& '1' & x"60";	-- LDA @352 	# Carrega o acumulador com o key 0
tmp(237) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador com o valor 0
tmp(238) := x"7" & "00" & '0' & '0' & x"E4";	-- JEQ %checa_limites_dezenas_de_milhares 	# Se for igual, vai para o label checa_limites_dezenas_de_milhares
tmp(239) := x"9" & "00" & '0' & '0' & x"F3";	-- JSR %adiciona_dezena_de_milhar 	# Se não for igual, vai para o label adiciona_dezena_de_milhar
tmp(240) := x"5" & "00" & '0'& '0' & x"2C";	-- STA @44 	# Armazena o valor do acumulador no endereço de Limite de dezenas de milhares
tmp(241) := x"6" & "00" & '0' & '0' & x"E0";	-- JMP %define_limites_dezenas_de_milhares 	# Se não for igual, volta para o label define_limites_dezenas_de_milhares
-- adiciona_dezena_de_milhar:
tmp(243) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(244) := x"1" & "00" & '0'& '0' & x"0F";	-- LDA @15 	# Carrega o acumulador com o endereço de Limite de dezena de milhar
tmp(245) := x"8" & "00" & '0'& '0' & x"34";	-- CEQ @52 	# Compara o valor do acumulador com o valor 9
tmp(246) := x"7" & "00"& '0' & '1' & x"00";	-- JEQ %limite_caso_20
tmp(247) := x"1" & "00" & '0'& '0' & x"2C";	-- LDA @44 	# Carrega o acumulador com o endereço de Limite de dezena de milhar
tmp(248) := x"8" & "00" & '0'& '0' & x"3B";	-- CEQ @59 	# Compara o valor do acumulador com o valor 9
tmp(249) := x"7" & "00" & '0' & '0' & x"FD";	-- JEQ %zera_dezena_de_milhar 	# Se for igual, vai para o label zera_dezena_de_milhar
tmp(250) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(251) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- zera_dezena_de_milhar:
tmp(253) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(254) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- limite_caso_20:
tmp(256) := x"1" & "00" & '0'& '0' & x"2C";	-- LDA @44 	# Carrega o acumulador com o endereço de Limite de dezena de milhar
tmp(257) := x"8" & "00" & '0'& '0' & x"35";	-- CEQ @53 	# Compara o valor do acumulador com o valor 9
tmp(258) := x"7" & "00" & '0' & '0' & x"FD";	-- JEQ %zera_dezena_de_milhar 	# Se for igual, vai para o label zera_dezena_de_milhar
tmp(259) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(260) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- define_limites_centenas_de_milhares:
tmp(262) := x"5" & "00" & '0'& '1' & x"FE";	-- STA @510 	# Limpando key 1
tmp(263) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(264) := x"5" & "00" & '0'& '1' & x"FD";	-- STA @509 	# Limpando key 0
tmp(265) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando key 0
tmp(266) := x"9" & "00" & '1' & '0' & x"6E";	-- JSR %atualiza_displays_limites 	# Vai para o label atualiza_displays_limites
-- checa_limites_centenas_de_milhares:
tmp(268) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(269) := x"5" & "00" & '0'& '1' & x"F8";	-- STA @504 	# liga o display unidade
tmp(270) := x"9" & "00" & '0' & '0' & x"47";	-- JSR %temporizador_1_segundo 	# Vai para o label temporizador_1_segundo
tmp(271) := x"1" & "00" & '0'& '0' & x"17";	-- LDA @23 	# Carrega o acumulador com o endereço de PISCA
tmp(272) := x"5" & "00" & '0'& '1' & x"F9";	-- STA @505 	# Desliga o display unidade
tmp(273) := x"1" & "00" & '0'& '1' & x"61";	-- LDA @353 	# Carrega o acumulador com o key 1
tmp(274) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(275) := x"7" & "00"& '0' & '1' & x"33";	-- JEQ %salva 	# Se for igual, vai para o label salva
tmp(276) := x"1" & "00" & '0'& '1' & x"62";	-- LDA @354 	# Carrega o acumulador com o key 2
tmp(277) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(278) := x"7" & "00"& '0' & '1' & x"41";	-- JEQ %salva_tempo 	# Se for igual, vai para o label salva
tmp(279) := x"1" & "00" & '0'& '1' & x"60";	-- LDA @352 	# Carrega o acumulador com o key 0
tmp(280) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador com o valor 0
tmp(281) := x"7" & "00"& '0' & '1' & x"0C";	-- JEQ %checa_limites_centenas_de_milhares 	# Se for igual, vai para o label checa_limites_centenas_de_milhares
tmp(282) := x"9" & "00"& '0' & '1' & x"1E";	-- JSR %adiciona_centena_de_milhar 	# Se não for igual, vai para o label adiciona_centena_de_milhar
tmp(283) := x"5" & "00" & '0'& '0' & x"2D";	-- STA @45 	# Armazena o valor do acumulador no endereço de Limite de centenas de milhares
tmp(284) := x"6" & "00"& '0' & '1' & x"06";	-- JMP %define_limites_centenas_de_milhares 	# Se não for igual, volta para o label define_limites_centenas_de_milhares
-- adiciona_centena_de_milhar:
tmp(286) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(287) := x"1" & "00" & '0'& '0' & x"2C";	-- LDA @44 	# Carrega o acumulador com o endereço de Limite de dezena de milhar
tmp(288) := x"8" & "00" & '0'& '0' & x"36";	-- CEQ @54 	# Compara o valor do acumulador com o valor 4
tmp(289) := x"C" & "00"& '0' & '1' & x"24";	-- JLT %limite_caso_24 	# Se for menor que 4, vai para o label limite_caso_24
tmp(290) := x"6" & "00"& '0' & '1' & x"2D";	-- JMP %especial_caso_24 	# Se não for menor que 4, vai para o label especial_caso_24
-- limite_caso_24:
tmp(292) := x"1" & "00" & '0'& '0' & x"2D";	-- LDA @45 	# Carrega o acumulador com o endereço de Limite de centena de milhar
tmp(293) := x"8" & "00" & '0'& '0' & x"34";	-- CEQ @52 	# Compara o valor do acumulador com o valor 2
tmp(294) := x"7" & "00"& '0' & '1' & x"2A";	-- JEQ %zera_centena_de_milhar 	# Se for igual, vai para o label zera_centena_de_milhar
tmp(295) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(296) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- zera_centena_de_milhar:
tmp(298) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 0 no acumulador
tmp(299) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- especial_caso_24:
tmp(301) := x"1" & "00" & '0'& '0' & x"2D";	-- LDA @45 	# Carrega o acumulador com o endereço de Limite de centena de milhar
tmp(302) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(303) := x"7" & "00"& '0' & '1' & x"2A";	-- JEQ %zera_centena_de_milhar 	# Se for igual, vai para o label zera_centena_de_milhar
tmp(304) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(305) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- salva:
tmp(307) := x"1" & "00" & '0'& '0' & x"2D";	-- LDA @45 	# Carrega o acumulador com o endereço de Limite de centena de milhar
tmp(308) := x"5" & "00" & '0'& '0' & x"0F";	-- STA @15 	# Armazena o valor do acumulador no endereço de Limite de dezena de milhar
tmp(309) := x"1" & "00" & '0'& '0' & x"2C";	-- LDA @44 	# Carrega o acumulador com o endereço de Limite de dezena de milhar
tmp(310) := x"5" & "00" & '0'& '0' & x"0E";	-- STA @14 	# Armazena o valor do acumulador no endereço de Limite de milhares
tmp(311) := x"1" & "00" & '0'& '0' & x"2B";	-- LDA @43 	# Carrega o acumulador com o endereço de Limite de milhares
tmp(312) := x"5" & "00" & '0'& '0' & x"0D";	-- STA @13 	# Armazena o valor do acumulador no endereço de Limite de centenas
tmp(313) := x"1" & "00" & '0'& '0' & x"2A";	-- LDA @42 	# Carrega o acumulador com o endereço de Limite de centenas
tmp(314) := x"5" & "00" & '0'& '0' & x"0C";	-- STA @12 	# Armazena o valor do acumulador no endereço de Limite de dezenas
tmp(315) := x"1" & "00" & '0'& '0' & x"29";	-- LDA @41 	# Carrega o acumulador com o endereço de Limite de dezenas
tmp(316) := x"5" & "00" & '0'& '0' & x"0B";	-- STA @11 	# Armazena o valor do acumulador no endereço de Limite de unidades
tmp(317) := x"1" & "00" & '0'& '0' & x"28";	-- LDA @40 	# Carrega o acumulador com o endereço de Limite de unidades
tmp(318) := x"5" & "00" & '0'& '0' & x"0A";	-- STA @10 	# Armazena o valor do acumulador no endereço de Limite de unidades
tmp(319) := x"6" & "00"& '0' & '1' & x"66";	-- JMP %reset_temp 	# Se não for igual, volta para o label define_limites_unidades
-- salva_tempo:
tmp(321) := x"1" & "00" & '0'& '0' & x"2D";	-- LDA @45 	# Carrega o acumulador com o endereço de Limite de centena de milhar
tmp(322) := x"5" & "00" & '0'& '0' & x"05";	-- STA @5 	# Armazena o valor do acumulador no endereço de Limite de dezena de milhar
tmp(323) := x"1" & "00" & '0'& '0' & x"2C";	-- LDA @44 	# Carrega o acumulador com o endereço de Limite de dezena de milhar
tmp(324) := x"5" & "00" & '0'& '0' & x"04";	-- STA @4 	# Armazena o valor do acumulador no endereço de Limite de milhares
tmp(325) := x"1" & "00" & '0'& '0' & x"2B";	-- LDA @43 	# Carrega o acumulador com o endereço de Limite de milhares
tmp(326) := x"5" & "00" & '0'& '0' & x"03";	-- STA @3 	# Armazena o valor do acumulador no endereço de Limite de centenas
tmp(327) := x"1" & "00" & '0'& '0' & x"2A";	-- LDA @42 	# Carrega o acumulador com o endereço de Limite de centenas
tmp(328) := x"5" & "00" & '0'& '0' & x"02";	-- STA @2 	# Armazena o valor do acumulador no endereço de Limite de dezenas
tmp(329) := x"1" & "00" & '0'& '0' & x"29";	-- LDA @41 	# Carrega o acumulador com o endereço de Limite de dezenas
tmp(330) := x"5" & "00" & '0'& '0' & x"01";	-- STA @1 	# Armazena o valor do acumulador no endereço de Limite de unidades
tmp(331) := x"1" & "00" & '0'& '0' & x"28";	-- LDA @40 	# Carrega o acumulador com o endereço de Limite de unidades
tmp(332) := x"5" & "00" & '0'& '0' & x"00";	-- STA @0 	# Armazena o valor do acumulador no endereço de Limite de unidades
tmp(333) := x"4" & "00" & '0'& '0' & x"55";	-- LDI $85 	# Carrega 85 no acumulador
tmp(334) := x"5" & "00" & '0'& '1' & x"00";	-- STA @256 	# Armazena o valor do acumulador nos LED 7 - 8
tmp(335) := x"1" & "00" & '0'& '1' & x"65";	-- LDA @357 	# Carrega o acumulador com o segundos
tmp(336) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(337) := x"7" & "00"& '0' & '1' & x"54";	-- JEQ %pre_salva_tempo_pt2
tmp(338) := x"6" & "00"& '0' & '1' & x"41";	-- JMP %salva_tempo
-- pre_salva_tempo_pt2:
tmp(340) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando key 0
-- salva_tempo_pt2:
tmp(342) := x"4" & "00" & '0'& '0' & x"55";	-- LDI $85 	# Carrega 85 no acumulador
tmp(343) := x"5" & "00" & '0'& '1' & x"00";	-- STA @256 	# Armazena o valor do acumulador nos LED 7 - 8
tmp(344) := x"1" & "00" & '0'& '1' & x"65";	-- LDA @357 	# Carrega o acumulador com o segundos
tmp(345) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(346) := x"7" & "00"& '0' & '1' & x"5D";	-- JEQ %pre_salva_tempo_pt3 	# Se não for igual, volta para o label define_limites_unidades
tmp(347) := x"6" & "00"& '0' & '1' & x"56";	-- JMP %salva_tempo_pt2
-- pre_salva_tempo_pt3:
tmp(349) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando key 0
-- salva_tempo_pt3:
tmp(351) := x"4" & "00" & '0'& '0' & x"AA";	-- LDI $170 	# Carrega 85 no acumulador
tmp(352) := x"5" & "00" & '0'& '1' & x"00";	-- STA @256 	# Armazena o valor do acumulador nos LED 7 - 8
tmp(353) := x"1" & "00" & '0'& '1' & x"65";	-- LDA @357 	# Carrega o acumulador com o segundos
tmp(354) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(355) := x"7" & "00"& '0' & '1' & x"66";	-- JEQ %reset_temp 	# Se não for igual, volta para o label define_limites_unidades
tmp(356) := x"6" & "00"& '0' & '1' & x"5F";	-- JMP %salva_tempo_pt3
-- reset_temp:
tmp(358) := x"1" & "00" & '0'& '0' & x"0A";	-- LDA @10 	# Carrega o acumulador com o endereço de Limite de unidades
tmp(359) := x"5" & "00" & '0'& '0' & x"28";	-- STA @40 	# Limpando endereço de temp 1
tmp(360) := x"1" & "00" & '0'& '0' & x"0C";	-- LDA @12 	# Carrega o acumulador com o endereço de Limite de CENTENAS
tmp(361) := x"5" & "00" & '0'& '0' & x"2A";	-- STA @42 	# Limpando endereço de temp 3
tmp(362) := x"1" & "00" & '0'& '0' & x"0B";	-- LDA @11 	# Carrega o acumulador com o endereço de Limite de CENTENAS
tmp(363) := x"5" & "00" & '0'& '0' & x"29";	-- STA @41 	# Limpando endereço de temp 2
tmp(364) := x"1" & "00" & '0'& '0' & x"0D";	-- LDA @13 	# Carrega o acumulador com o endereço de Limite de CENTENAS
tmp(365) := x"5" & "00" & '0'& '0' & x"2B";	-- STA @43 	# Limpando endereço de temp 4
tmp(366) := x"1" & "00" & '0'& '0' & x"0E";	-- LDA @14 	# Carrega o acumulador com o endereço de Limite de CENTENAS
tmp(367) := x"5" & "00" & '0'& '0' & x"2C";	-- STA @44 	# Limpando endereço de temp 5
tmp(368) := x"1" & "00" & '0'& '0' & x"0F";	-- LDA @15 	# Carrega o acumulador com o endereço de Limite de CENTENAS
tmp(369) := x"5" & "00" & '0'& '0' & x"2D";	-- STA @45 	# Limpando endereço de temp 6
tmp(370) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 85 no acumulador
tmp(371) := x"5" & "00" & '0'& '1' & x"00";	-- STA @256 	# Armazena o valor do acumulador nos LED 7 - 8
tmp(372) := x"6" & "00"& '0' & '1' & x"76";	-- JMP %pre_le_key
-- pre_le_key:
tmp(374) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(375) := x"5" & "00" & '0'& '1' & x"FE";	-- STA @510 	# Limpando key 1
tmp(376) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega 1 no acumulador
tmp(377) := x"5" & "00" & '0'& '1' & x"F9";	-- STA @505 	# Liga o display 0
tmp(378) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays
tmp(379) := x"6" & "00"& '0' & '1' & x"7D";	-- JMP %le_key 	# Vai para o label le_key
-- le_key:
tmp(381) := x"1" & "00" & '0'& '1' & x"65";	-- LDA @357 	# Carrega o acumulador com o segundos
tmp(382) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(383) := x"7" & "00"& '0' & '1' & x"A0";	-- JEQ %incrementa_unidade 	# Se for igual, vai para o label incrementa
tmp(384) := x"1" & "00" & '0'& '1' & x"61";	-- LDA @353 	# Carrega o acumulador com o key 1
tmp(385) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(386) := x"7" & "00" & '0' & '0' & x"6D";	-- JEQ %define_limites_unidades 	# Se for igual, vai para o label incrementa
tmp(387) := x"9" & "00"& '0' & '1' & x"8A";	-- JSR %checa_op 	# checa se é + ou -
tmp(388) := x"9" & "00"& '0' & '1' & x"95";	-- JSR %checa_timer 	# checa se ta ligado ou nao
tmp(389) := x"1" & "00" & '0'& '1' & x"64";	-- LDA @356		# Carrega o acumulador com o endereço de fpga_reset
tmp(390) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(391) := x"7" & "00" & '1' & '0' & x"9F";	-- JEQ %RESET_FPGA 	# Se for igual, vai para o label RESET_FPGA
tmp(392) := x"6" & "00"& '0' & '1' & x"7D";	-- JMP %le_key 	# Se não for igual, volta para o label le_key
-- checa_op:
tmp(394) := x"1" & "00" & '0'& '1' & x"42";	-- LDA @322 	# Carrega o acumulador com o endereço de SW9
tmp(395) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador com o valor 0
tmp(396) := x"7" & "00"& '0' & '1' & x"91";	-- JEQ %mais 	# Se for igual, vai para o label le_key
tmp(397) := x"4" & "00" & '0'& '0' & x"01";	-- LDI $1 	# Carrega o acumulador com o valor 1
tmp(398) := x"5" & "00" & '0'& '1' & x"02";	-- STA @258 	# Liga led 9
tmp(399) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- mais:
tmp(401) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega o acumulador com o valor 1
tmp(402) := x"5" & "00" & '0'& '1' & x"02";	-- STA @258 	# Liga led 9
tmp(403) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- checa_timer:
tmp(405) := x"1" & "00" & '0'& '1' & x"41";	-- LDA @321 	# Carrega o acumulador com o endereço de SW8
tmp(406) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador com o valor 0
tmp(407) := x"7" & "00"& '0' & '1' & x"9C";	-- JEQ %desativado 	# Se for igual, vai para o label desativado
tmp(408) := x"4" & "00" & '0'& '0' & x"01";	-- LDI $1 	# Carrega o acumulador com o valor 1
tmp(409) := x"5" & "00" & '0'& '1' & x"01";	-- STA @257 	# Liga led 8
tmp(410) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- desativado:
tmp(412) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega o acumulador com o valor 1
tmp(413) := x"5" & "00" & '0'& '1' & x"01";	-- STA @257 	# Liga led 8
tmp(414) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- incrementa_unidade:
tmp(416) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando key 0
tmp(417) := x"1" & "00" & '0'& '1' & x"42";	-- LDA @322 	# Carrega o acumulador com o endereço de SW9
tmp(418) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(419) := x"7" & "00"& '0' & '1' & x"AD";	-- JEQ %sub_unidade 	# Se for igual, vai para o label sub_unidade
tmp(420) := x"1" & "00" & '0'& '0' & x"00";	-- LDA @0 	# Carrega o acumulador com o endereço de unidade
tmp(421) := x"8" & "00" & '0'& '0' & x"3B";	-- CEQ @59 	# Compara o valor do acumulador com o valor 9
tmp(422) := x"7" & "00"& '0' & '1' & x"B4";	-- JEQ %incrementa_dezena 	# Se for igual, vai para o label incrementa_dezena
tmp(423) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(424) := x"5" & "00" & '0'& '0' & x"00";	-- STA @0 	# Armazena o valor do acumulador no endereço de unidade
tmp(425) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carrega o acumulador com o valor 1
tmp(426) := x"5" & "00" & '0'& '1' & x"02";	-- STA @258 	# Desliga led 9
tmp(427) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, vai para o label atualiza_unidade
-- sub_unidade:
tmp(429) := x"1" & "00" & '0'& '0' & x"00";	-- LDA @0 	# Carrega o acumulador com o endereço de unidade
tmp(430) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador com o valor 0
tmp(431) := x"7" & "00"& '0' & '1' & x"BE";	-- JEQ %decremeta_dezena 	# Se for igual, vai para o label decremeta_dezena
tmp(432) := x"3" & "00" & '0'& '0' & x"33";	-- SUB @51 	# Subtrai 1 no acumulador
tmp(433) := x"5" & "00" & '0'& '0' & x"00";	-- STA @0 	# Armazena o valor do acumulador no endereço de unidade
tmp(434) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, vai para o label atualiza_unidade
-- incrementa_dezena:
tmp(436) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0
tmp(437) := x"5" & "00" & '0'& '0' & x"00";	-- STA @0 	# Limpando endereço de unidade
tmp(438) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando Key 0
tmp(439) := x"1" & "00" & '0'& '0' & x"01";	-- LDA @1 	# Carregar o acumulador com o endereço da dezena
tmp(440) := x"8" & "00" & '0'& '0' & x"37";	-- CEQ @55 	# Compara o valor do acumulador (dezena) com o valor 9
tmp(441) := x"7" & "00"& '0' & '1' & x"C8";	-- JEQ %incrementa_centena 	# Se for igual a 9, vai para o incrementa_centena
tmp(442) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(443) := x"5" & "00" & '0'& '0' & x"01";	-- STA @1 	# Armazena o valor do acumulador no endereço das dezenas
tmp(444) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, volta para o label atualiza_displays
-- decremeta_dezena:
tmp(446) := x"4" & "00" & '0'& '0' & x"09";	-- LDI $9
tmp(447) := x"5" & "00" & '0'& '0' & x"00";	-- STA @0 	# Limpando endereço de unidade
tmp(448) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando Key 0
tmp(449) := x"1" & "00" & '0'& '0' & x"01";	-- LDA @1 	# Carregar o acumulador com o endereço da dezena
tmp(450) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador (dezena) com o valor 0
tmp(451) := x"7" & "00"& '0' & '1' & x"D2";	-- JEQ %decremeta_centena 	# Se for igual a 0, vai para o decremeta_centena
tmp(452) := x"3" & "00" & '0'& '0' & x"33";	-- SUB @51 	# Subtrai 1 no acumulador
tmp(453) := x"5" & "00" & '0'& '0' & x"01";	-- STA @1 	# Armazena o valor do acumulador no endereço das dezenas
tmp(454) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, volta para o label atualiza_displays
-- incrementa_centena:
tmp(456) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0
tmp(457) := x"5" & "00" & '0'& '0' & x"01";	-- STA @1 	# Limpando endereço de dezena
tmp(458) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando Key 0
tmp(459) := x"1" & "00" & '0'& '0' & x"02";	-- LDA @2 	# Carregar o acumulador com o endereço da centena
tmp(460) := x"8" & "00" & '0'& '0' & x"3B";	-- CEQ @59 	# Compara o valor do acumulador (centena) com o valor 9
tmp(461) := x"7" & "00"& '0' & '1' & x"DC";	-- JEQ %incrementa_milhar 	# Se for igual a 9, vai para o incrementa_milhar
tmp(462) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(463) := x"5" & "00" & '0'& '0' & x"02";	-- STA @2 	# Armazena o valor do acumulador no endereço das centenas
tmp(464) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, volta para o label atualiza_displays
-- decremeta_centena:
tmp(466) := x"4" & "00" & '0'& '0' & x"05";	-- LDI $5
tmp(467) := x"5" & "00" & '0'& '0' & x"01";	-- STA @1 	# Limpando endereço de dezena
tmp(468) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando Key 0
tmp(469) := x"1" & "00" & '0'& '0' & x"02";	-- LDA @2 	# Carregar o acumulador com o endereço da centena
tmp(470) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador (centena) com o valor 0
tmp(471) := x"7" & "00"& '0' & '1' & x"E6";	-- JEQ %decremeta_milhar 	# Se for igual a 0, vai para o decremeta_milhar
tmp(472) := x"3" & "00" & '0'& '0' & x"33";	-- SUB @51 	# Subtrai 1 no acumulador
tmp(473) := x"5" & "00" & '0'& '0' & x"02";	-- STA @2 	# Armazena o valor do acumulador no endereço das centenas
tmp(474) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, volta para o label atualiza_displays
-- incrementa_milhar:
tmp(476) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0
tmp(477) := x"5" & "00" & '0'& '0' & x"02";	-- STA @2 	# Limpando endereço de centena
tmp(478) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando Key 0
tmp(479) := x"1" & "00" & '0'& '0' & x"03";	-- LDA @3 	# Carregar o acumulador com o endereço da milhares
tmp(480) := x"8" & "00" & '0'& '0' & x"37";	-- CEQ @55 	# Compara o valor do acumulador (dezena) com o valor 9
tmp(481) := x"7" & "00"& '0' & '1' & x"F0";	-- JEQ %incrementa_dezena_de_milhar 	# Se for igual a 9, vai para o incrementa_dezena_de_milhar
tmp(482) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(483) := x"5" & "00" & '0'& '0' & x"03";	-- STA @3 	# Armazena o valor do acumulador no endereço das milhares
tmp(484) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, volta para o label atualiza_unidade
-- decremeta_milhar:
tmp(486) := x"4" & "00" & '0'& '0' & x"09";	-- LDI $9
tmp(487) := x"5" & "00" & '0'& '0' & x"02";	-- STA @2 	# Limpando endereço de centena
tmp(488) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando Key 0
tmp(489) := x"1" & "00" & '0'& '0' & x"03";	-- LDA @3 	# Carregar o acumulador com o endereço da milhares
tmp(490) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador (dezena) com o valor 0
tmp(491) := x"7" & "00" & '1' & '0' & x"03";	-- JEQ %decremeta_dezena_de_milhar 	# Se for igual a 0, vai para o decremeta_dezena_de_milhar
tmp(492) := x"3" & "00" & '0'& '0' & x"33";	-- SUB @51 	# Subtrai 1 no acumulador
tmp(493) := x"5" & "00" & '0'& '0' & x"03";	-- STA @3 	# Armazena o valor do acumulador no endereço das milhares
tmp(494) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, volta para o label atualiza_unidade
-- incrementa_dezena_de_milhar:
tmp(496) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0
tmp(497) := x"5" & "00" & '0'& '0' & x"03";	-- STA @3 	# Limpando endereço de milhar (RAM 3)
tmp(498) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando Key 0
tmp(499) := x"1" & "00" & '0'& '0' & x"05";	-- LDA @5 	# Carregar o acumulador com o endereço da centena de milhar
tmp(500) := x"8" & "00" & '0'& '0' & x"34";	-- CEQ @52 	# Compara o valor do acumulador (dezena) com o valor 2
tmp(501) := x"7" & "00"& '0' & '1' & x"FE";	-- JEQ %outro_incremente_dezena_de_milhar 	# Se for igual a 2, vai para o incremenoutro_incremente_dezena_de_milharta_centena_milhar
tmp(502) := x"1" & "00" & '0'& '0' & x"04";	-- LDA @4 	# Carregar o acumulador com o endereço da dezena de milhar
tmp(503) := x"8" & "00" & '0'& '0' & x"3B";	-- CEQ @59 	# Compara o valor do acumulador (dezena) com o valor 9
tmp(504) := x"7" & "00" & '1' & '0' & x"0D";	-- JEQ %incrementa_centena_milhar 	# Se for igual a 9, vai para o incrementa_centena_milhar
-- volta:
tmp(506) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(507) := x"5" & "00" & '0'& '0' & x"04";	-- STA @4 	# Armazena o valor do acumulador no endereço das milhares
tmp(508) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, volta para o label atualiza_displays
-- outro_incremente_dezena_de_milhar:
tmp(510) := x"1" & "00" & '0'& '0' & x"04";	-- LDA @4 	# Carregar o acumulador com o endereço da dezena de milhar
tmp(511) := x"8" & "00" & '0'& '0' & x"35";	-- CEQ @53 	# Compara o valor do acumulador (dezena) com o valor 9
tmp(512) := x"7" & "00" & '1' & '0' & x"0D";	-- JEQ %incrementa_centena_milhar 	# Se for igual a 9, vai para o incrementa_centena_milhar
tmp(513) := x"6" & "00"& '0' & '1' & x"FA";	-- JMP %volta 	# Se não for igual, volta para o label volta
-- decremeta_dezena_de_milhar:
tmp(515) := x"4" & "00" & '0'& '0' & x"05";	-- LDI $5
tmp(516) := x"5" & "00" & '0'& '0' & x"03";	-- STA @3 	# Limpando endereço de milhar (RAM 3)
tmp(517) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando Key 0
tmp(518) := x"1" & "00" & '0'& '0' & x"04";	-- LDA @4 	# Carregar o acumulador com o endereço da dezena de milhar
tmp(519) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador (dezena) com o valor 0
tmp(520) := x"7" & "00" & '1' & '0' & x"17";	-- JEQ %decremeta_centena_milhar 	# Se for igual a 0, vai para o decremeta_centena_milhar
tmp(521) := x"3" & "00" & '0'& '0' & x"33";	-- SUB @51 	# Subtrai 1 no acumulador
tmp(522) := x"5" & "00" & '0'& '0' & x"04";	-- STA @4 	# Armazena o valor do acumulador no endereço das milhares
tmp(523) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, volta para o label atualiza_displays
-- incrementa_centena_milhar:
tmp(525) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0
tmp(526) := x"5" & "00" & '0'& '0' & x"04";	-- STA @4 	# Limpando endereço de dezena de milhar
tmp(527) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando Key 0
tmp(528) := x"1" & "00" & '0'& '0' & x"05";	-- LDA @5 	# Carregar o acumulador com o endereço da centena
tmp(529) := x"8" & "00" & '0'& '0' & x"34";	-- CEQ @52 	# Compara o valor do acumulador (centena) com o valor 9
tmp(530) := x"7" & "00" & '1' & '0' & x"29";	-- JEQ %zerou 	# Se for igual a 9, vai para o atualiza_displays
tmp(531) := x"2" & "00" & '0'& '0' & x"33";	-- SOMA @51 	# Soma 1 no acumulador
tmp(532) := x"5" & "00" & '0'& '0' & x"05";	-- STA @5 	# Armazena o valor do acumulador no endereço das centenas
tmp(533) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, volta para o label atualiza_displays
-- decremeta_centena_milhar:
tmp(535) := x"1" & "00" & '0'& '0' & x"05";	-- LDA @5 	# Carrega o acumulador com o endereço de centena de milhar
tmp(536) := x"8" & "00" & '0'& '0' & x"34";	-- CEQ @52 	# Compara o valor do acumulador com o valor 2 (limite de centena de milhar)
tmp(537) := x"7" & "00" & '1' & '0' & x"25";	-- JEQ %caso20 	# Se for igual, vai para o label caso20
tmp(538) := x"4" & "00" & '0'& '0' & x"03";	-- LDI $3
tmp(539) := x"5" & "00" & '0'& '0' & x"04";	-- STA @4 	# Limpando endereço de dezena de milhar
-- volta_caso20:
tmp(541) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando Key 0
tmp(542) := x"1" & "00" & '0'& '0' & x"05";	-- LDA @5 	# Carregar o acumulador com o endereço da centena
tmp(543) := x"8" & "00" & '0'& '0' & x"32";	-- CEQ @50 	# Compara o valor do acumulador (centena) com o valor 0
tmp(544) := x"7" & "00" & '1' & '0' & x"29";	-- JEQ %zerou 	# Se for igual a 0, vai para o atualiza_displays
tmp(545) := x"3" & "00" & '0'& '0' & x"33";	-- SUB @51 	# Subtrai 1 no acumulador
tmp(546) := x"5" & "00" & '0'& '0' & x"05";	-- STA @5 	# Armazena o valor do acumulador no endereço das centenas
tmp(547) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Se não for igual, volta para o label atualiza_displays
-- caso20:
tmp(549) := x"4" & "00" & '0'& '0' & x"09";	-- LDI $9  
tmp(550) := x"5" & "00" & '0'& '0' & x"04";	-- STA @4 	# Limpando endereço de dezena de milhar
tmp(551) := x"6" & "00" & '1' & '0' & x"1D";	-- JMP %volta_caso20 	# Se não for igual, volta para o label volta_caso20
-- zerou:
tmp(553) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0
tmp(554) := x"5" & "00" & '0'& '0' & x"05";	-- STA @5 	# Limpando endereço de centena de milhar
tmp(555) := x"5" & "00" & '0'& '0' & x"04";	-- STA @4 	# Limpando endereço de dezena de milhar
tmp(556) := x"5" & "00" & '0'& '0' & x"03";	-- STA @3 	# Limpando endereço de milhar
tmp(557) := x"5" & "00" & '0'& '0' & x"02";	-- STA @2 	# Limpando endereço de centena
tmp(558) := x"5" & "00" & '0'& '0' & x"01";	-- STA @1 	# Limpando endereço de dezena
tmp(559) := x"5" & "00" & '0'& '0' & x"00";	-- STA @0 	# Limpando endereço de unidade
tmp(560) := x"1" & "00" & '0'& '1' & x"42";	-- LDA @322 	# Carrega o acumulador com o endereço de SW9
tmp(561) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(562) := x"7" & "00" & '1' & '0' & x"AB";	-- JEQ %final 	# Se for igual, vai para o label final
tmp(563) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando Key 0
tmp(564) := x"5" & "00" & '0'& '1' & x"FE";	-- STA @510 	# Limpando Key 1
tmp(565) := x"4" & "00" & '0'& '0' & x"01";	-- LDI $1 	# Carrega 2 no acumulador
tmp(566) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Vai para o label atualiza_displays
-- atualiza_displays:
tmp(568) := x"1" & "00" & '0'& '0' & x"00";	-- LDA @0 	# Carrega o acumulador com o endereço de unidade
tmp(569) := x"5" & "00" & '0'& '1' & x"20";	-- STA @288 	# Armazena o valor do acumulador no endereço do HEX0
tmp(570) := x"1" & "00" & '0'& '0' & x"01";	-- LDA @1 	# Carrega o acumulador com o endereço de dezena
tmp(571) := x"5" & "00" & '0'& '1' & x"21";	-- STA @289 	# Armazena o valor do acumulador no endereço do HEX1
tmp(572) := x"1" & "00" & '0'& '0' & x"02";	-- LDA @2 	# Carrega o acumulador com o endereço de centena
tmp(573) := x"5" & "00" & '0'& '1' & x"22";	-- STA @290 	# Armazena o valor do acumulador no endereço do HEX2
tmp(574) := x"1" & "00" & '0'& '0' & x"03";	-- LDA @3 	# Carrega o acumulador com o endereço de milhar
tmp(575) := x"5" & "00" & '0'& '1' & x"23";	-- STA @291 	# Armazena o valor do acumulador no endereço do HEX3
tmp(576) := x"1" & "00" & '0'& '0' & x"04";	-- LDA @4 	# Carrega o acumulador com o endereço de dezena de milhar
tmp(577) := x"5" & "00" & '0'& '1' & x"24";	-- STA @292 	# Armazena o valor do acumulador no endereço do HEX4
tmp(578) := x"1" & "00" & '0'& '0' & x"05";	-- LDA @5 	# Carrega o acumulador com o endereço de centena de milhar
tmp(579) := x"5" & "00" & '0'& '1' & x"25";	-- STA @293 	# Armazena o valor do acumulador no endereço do HEX5
tmp(580) := x"9" & "00" & '1' & '0' & x"48";	-- JSR %atualiza_vga 	# Vai para o label atualiza_vga
tmp(581) := x"9" & "00" & '1' & '0' & x"7C";	-- JSR %verifica_centena_de_milhar 	# Vai para o label verifica_centena_de_milhar
tmp(582) := x"6" & "00"& '0' & '1' & x"7D";	-- JMP %le_key 	# Vai para o label le_key
-- atualiza_vga:
tmp(584) := x"4" & "00" & '0'& '0' & x"10";	-- LDI $16 	# Carrega o acumulador com o valor 16
tmp(585) := x"2" & "00" & '0'& '0' & x"00";	-- SOMA @0 	# Soma 16 no acumulador
tmp(586) := x"5" & "00" & '0'& '0' & x"82";	-- STA @ 130 	# Armazena o valor do acumulador no endereço dos caracteres
tmp(587) := x"4" & "00" & '0'& '0' & x"0D";	-- LDI $13 	# Carrega o acumulador com o valor 13
tmp(588) := x"5" & "00" & '0'& '0' & x"81";	-- STA @129 	# Armazena o valor do acumulador na COLUNA
tmp(589) := x"5" & "00" & '0'& '0' & x"83";	-- STA @131 	# HABILITA VGA
tmp(590) := x"4" & "00" & '0'& '0' & x"10";	-- LDI $16 	# Carrega o acumulador com o valor 16
tmp(591) := x"2" & "00" & '0'& '0' & x"01";	-- SOMA @1 	# Soma 16 no acumulador
tmp(592) := x"5" & "00" & '0'& '0' & x"82";	-- STA @ 130 	# Armazena o valor do acumulador no endereço dos caracteres
tmp(593) := x"4" & "00" & '0'& '0' & x"0C";	-- LDI $12 	# Carrega o acumulador com o valor 12
tmp(594) := x"5" & "00" & '0'& '0' & x"81";	-- STA @129 	# Armazena o valor do acumulador na COLUNA
tmp(595) := x"5" & "00" & '0'& '0' & x"83";	-- STA @131 	# HABILITA VGA
tmp(596) := x"4" & "00" & '0'& '0' & x"10";	-- LDI $16 	# Carrega o acumulador com o valor 16
tmp(597) := x"2" & "00" & '0'& '0' & x"02";	-- SOMA @2 	# Soma 16 no acumulador
tmp(598) := x"5" & "00" & '0'& '0' & x"82";	-- STA @ 130 	# Armazena o valor do acumulador no endereço dos caracteres
tmp(599) := x"4" & "00" & '0'& '0' & x"0A";	-- LDI $10 	# Carrega o acumulador com o valor 12
tmp(600) := x"5" & "00" & '0'& '0' & x"81";	-- STA @129 	# Armazena o valor do acumulador na COLUNA
tmp(601) := x"5" & "00" & '0'& '0' & x"83";	-- STA @131 	# HABILITA VGA
tmp(602) := x"4" & "00" & '0'& '0' & x"10";	-- LDI $16 	# Carrega o acumulador com o valor 16
tmp(603) := x"2" & "00" & '0'& '0' & x"03";	-- SOMA @3 	# Soma 16 no acumulador
tmp(604) := x"5" & "00" & '0'& '0' & x"82";	-- STA @ 130 	# Armazena o valor do acumulador no endereço dos caracteres
tmp(605) := x"4" & "00" & '0'& '0' & x"09";	-- LDI $9 	# Carrega o acumulador com o valor 12
tmp(606) := x"5" & "00" & '0'& '0' & x"81";	-- STA @129 	# Armazena o valor do acumulador na COLUNA
tmp(607) := x"5" & "00" & '0'& '0' & x"83";	-- STA @131 	# HABILITA VGA
tmp(608) := x"4" & "00" & '0'& '0' & x"10";	-- LDI $16 	# Carrega o acumulador com o valor 16
tmp(609) := x"2" & "00" & '0'& '0' & x"04";	-- SOMA @4 	# Soma 16 no acumulador
tmp(610) := x"5" & "00" & '0'& '0' & x"82";	-- STA @ 130 	# Armazena o valor do acumulador no endereço dos caracteres
tmp(611) := x"4" & "00" & '0'& '0' & x"07";	-- LDI $7 	# Carrega o acumulador com o valor 12
tmp(612) := x"5" & "00" & '0'& '0' & x"81";	-- STA @129 	# Armazena o valor do acumulador na COLUNA
tmp(613) := x"5" & "00" & '0'& '0' & x"83";	-- STA @131 	# HABILITA VGA
tmp(614) := x"4" & "00" & '0'& '0' & x"10";	-- LDI $16 	# Carrega o acumulador com o valor 16
tmp(615) := x"2" & "00" & '0'& '0' & x"05";	-- SOMA @5 	# Soma 16 no acumulador
tmp(616) := x"5" & "00" & '0'& '0' & x"82";	-- STA @ 130 	# Armazena o valor do acumulador no endereço dos caracteres
tmp(617) := x"4" & "00" & '0'& '0' & x"06";	-- LDI $6 	# Carrega o acumulador com o valor 12
tmp(618) := x"5" & "00" & '0'& '0' & x"81";	-- STA @129 	# Armazena o valor do acumulador na COLUNA
tmp(619) := x"5" & "00" & '0'& '0' & x"83";	-- STA @131 	# HABILITA VGA
tmp(620) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- atualiza_displays_limites:
tmp(622) := x"1" & "00" & '0'& '0' & x"28";	-- LDA @40 	# Carrega o acumulador com o Limites das unidades
tmp(623) := x"5" & "00" & '0'& '1' & x"20";	-- STA @288 	# Armazena o valor do acumulador no endereço do HEX0
tmp(624) := x"1" & "00" & '0'& '0' & x"29";	-- LDA @41 	# Carrega o acumulador com o Limites das dezenas
tmp(625) := x"5" & "00" & '0'& '1' & x"21";	-- STA @289 	# Armazena o valor do acumulador no endereço do HEX1
tmp(626) := x"1" & "00" & '0'& '0' & x"2A";	-- LDA @42 	# Carrega o acumulador com o Limites de centena
tmp(627) := x"5" & "00" & '0'& '1' & x"22";	-- STA @290 	# Armazena o valor do acumulador no endereço do HEX2
tmp(628) := x"1" & "00" & '0'& '0' & x"2B";	-- LDA @43 	# Carrega o acumulador com o Limites de milhar
tmp(629) := x"5" & "00" & '0'& '1' & x"23";	-- STA @291 	# Armazena o valor do acumulador no endereço do HEX3
tmp(630) := x"1" & "00" & '0'& '0' & x"2C";	-- LDA @44 	# Carrega o acumulador com o Limites de dezena de milhar
tmp(631) := x"5" & "00" & '0'& '1' & x"24";	-- STA @292 	# Armazena o valor do acumulador no endereço do HEX4
tmp(632) := x"1" & "00" & '0'& '0' & x"2D";	-- LDA @45 	# Carrega o acumulador com o Limites de centena de milhar
tmp(633) := x"5" & "00" & '0'& '1' & x"25";	-- STA @293 	# Armazena o valor do acumulador no endereço do HEX5
tmp(634) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- verifica_centena_de_milhar:
tmp(636) := x"1" & "00" & '0'& '1' & x"41";	-- LDA @321 	# Carrega o acumulador com o endereço de SW8
tmp(637) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 0
tmp(638) := x"7" & "00" & '1' & '0' & x"81";	-- JEQ %continua_verifica_centena_de_milhar 	# Se for igual, vai para o label continua_verifica_centena_de_milhar
tmp(639) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- continua_verifica_centena_de_milhar: 
tmp(641) := x"1" & "00" & '0'& '0' & x"05";	-- LDA @5 	# Carrega o acumulador com o endereço de centena de milhar
tmp(642) := x"8" & "00" & '0'& '0' & x"0F";	-- CEQ @15 	# Compara o valor do acumulador com o valor maximo de centena de milhar
tmp(643) := x"7" & "00" & '1' & '0' & x"86";	-- JEQ %verifica_dezena_de_milhar 	# Se for igual, vai para o label verifica_dezena_de_milhar
tmp(644) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- verifica_dezena_de_milhar:
tmp(646) := x"1" & "00" & '0'& '0' & x"04";	-- LDA @4 	# Carrega o acumulador com o endereço de dezena de milhar
tmp(647) := x"8" & "00" & '0'& '0' & x"0E";	-- CEQ @14 	# Compara o valor do acumulador com o valor maximo de dezena de milhar
tmp(648) := x"7" & "00" & '1' & '0' & x"8B";	-- JEQ %verifica_milhar 	# Se for igual, vai para o label verifica_milhar
tmp(649) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- verifica_milhar:
tmp(651) := x"1" & "00" & '0'& '0' & x"03";	-- LDA @3 	# Carrega o acumulador com o endereço de milhar
tmp(652) := x"8" & "00" & '0'& '0' & x"0D";	-- CEQ @13 	# Compara o valor do acumulador com o valor maximo de milhar
tmp(653) := x"7" & "00" & '1' & '0' & x"90";	-- JEQ %verifica_centena 	# Se for igual, vai para o label verifica_centena
tmp(654) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- verifica_centena:
tmp(656) := x"1" & "00" & '0'& '0' & x"02";	-- LDA @2 	# Carrega o acumulador com o endereço de centena
tmp(657) := x"8" & "00" & '0'& '0' & x"0C";	-- CEQ @12 	# Compara o valor do acumulador com o valor maximo de centena
tmp(658) := x"7" & "00" & '1' & '0' & x"95";	-- JEQ %verifica_dezena 	# Se for igual, vai para o label verifica_dezena
tmp(659) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- verifica_dezena:
tmp(661) := x"1" & "00" & '0'& '0' & x"01";	-- LDA @1 	# Carrega o acumulador com o endereço de dezena
tmp(662) := x"8" & "00" & '0'& '0' & x"0B";	-- CEQ @11 	# Compara o valor do acumulador com o valor maximo de dezena
tmp(663) := x"7" & "00" & '1' & '0' & x"9A";	-- JEQ %verifica_unidade 	# Se for igual, vai para o label verifica_unidade
tmp(664) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- verifica_unidade:
tmp(666) := x"1" & "00" & '0'& '0' & x"00";	-- LDA @0 	# Carrega o acumulador com o endereço de unidade
tmp(667) := x"8" & "00" & '0'& '0' & x"0A";	-- CEQ @10 	# Compara o valor do acumulador com o valor maximo de unidade
tmp(668) := x"7" & "00" & '1' & '0' & x"AB";	-- JEQ %final 	# Se for igual, vai para o label final
tmp(669) := x"A" & "00" & '0' & '0' & x"00";	-- RET
-- RESET_FPGA:
tmp(671) := x"5" & "00" & '0'& '1' & x"FF";	-- STA @511 	# Limpando key 0
tmp(672) := x"5" & "00" & '0'& '1' & x"FE";	-- STA @510 	# Limpando key 1
tmp(673) := x"5" & "00" & '0'& '1' & x"FC";	-- STA @508 	# Limpando reset_key
tmp(674) := x"4" & "00" & '0'& '0' & x"00";	-- LDI $0 	# Carregando 0 no acumulador
tmp(675) := x"5" & "00" & '0'& '1' & x"02";	-- STA @258 	# Desliga led 9
tmp(676) := x"5" & "00" & '0'& '1' & x"01";	-- STA @257 	# Desliga o led 8
tmp(677) := x"5" & "00" & '0'& '1' & x"00";	-- STA @256 	# Desliga o led 7 ao led 0
tmp(678) := x"5" & "00" & '1' & '1' & x"FF";	-- STA @1023 	# Desliga o BUZZER
tmp(679) := x"4" & "00" & '0'& '0' & x"07";	-- LDI $7 	# Carregando 7 no acumulador
tmp(680) := x"5" & "00" & '0'& '0' & x"84";	-- STA @132 	# Carregando 7 na COR
tmp(681) := x"6" & "00" & '1' & '0' & x"38";	-- JMP %atualiza_displays 	# Vai para o label atualiza_displays
-- final:
tmp(683) := x"4" & "00" & '0'& '0' & x"01";	-- LDI $1 	# Carrega 2 no acumulador
tmp(684) := x"5" & "00" & '0'& '0' & x"84";	-- STA @132 	# Carrega 2 na COR
tmp(685) := x"9" & "00" & '1' & '0' & x"48";	-- JSR %atualiza_vga 	# Vai para o label atualiza_vga
tmp(686) := x"4" & "00" & '0'& '0' & x"01";	-- LDI $1 	# Carrega 1 no acumulador
tmp(687) := x"5" & "00" & '1' & '1' & x"FF";	-- STA @1023 	# Liga o BUZZER
tmp(688) := x"1" & "00" & '0'& '0' & x"33";	-- LDA @51 	# Carrega 1 no acumulador
tmp(689) := x"5" & "00" & '0'& '1' & x"02";	-- STA @258 	# Liga led 9
tmp(690) := x"5" & "00" & '0'& '1' & x"01";	-- STA @257 	# Liga o led 8
tmp(691) := x"4" & "00" & '0'& '0' & x"FF";	-- LDI $255 	# Carrega 255 no acumulador
tmp(692) := x"5" & "00" & '0'& '1' & x"00";	-- STA @256 	# Liga o led 7 ao led 0
tmp(693) := x"1" & "00" & '0'& '1' & x"64";	-- LDA @356		# Carrega o acumulador com o endereço de fpga_reset
tmp(694) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(695) := x"7" & "00" & '1' & '0' & x"9F";	-- JEQ %RESET_FPGA 	# Se for igual, vai para o label RESET_FPGA
tmp(696) := x"1" & "00" & '0'& '1' & x"61";	-- LDA @353 	# Carrega o acumulador com o key 1
tmp(697) := x"8" & "00" & '0'& '0' & x"33";	-- CEQ @51 	# Compara o valor do acumulador com o valor 1
tmp(698) := x"7" & "00" & '0' & '0' & x"6D";	-- JEQ %define_limites_unidades 	# Se for igual, vai para o label incrementa
tmp(699) := x"6" & "00"& '0' & '1' & x"7D";	-- JMP %le_key 	# Se não for igual, volta para o label le_key

        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;